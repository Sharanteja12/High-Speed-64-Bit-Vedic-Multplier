module csa_64 (a,b,c,s,cout);

input [63:0]a,b,c;
output [64:0] s;
output cout ;

wire [63:0] s1,c1;
fa e1(a[0],b[0],c[0],s1[0],c1[0]);
fa e2(a[1],b[1],c[1],s1[1],c1[1]);
fa e3(a[2],b[2],c[2],s1[2],c1[2]);
fa e4(a[3],b[3],c[3],s1[3],c1[3]);
fa e5(a[4],b[4],c[4],s1[4],c1[4]);
fa e6(a[5],b[5],c[5],s1[5],c1[5]);
fa e7(a[6],b[6],c[6],s1[6],c1[6]);
fa e8(a[7],b[7],c[7],s1[7],c1[7]);

fa e9(a[8],b[8],c[8],s1[8],c1[8]);
fa e10(a[9],b[9],c[9],s1[9],c1[9]);
fa e11(a[10],b[10],c[10],s1[10],c1[10]);
fa e12(a[11],b[11],c[11],s1[11],c1[11]);
fa e13(a[12],b[12],c[12],s1[12],c1[12]);
fa e14(a[13],b[13],c[13],s1[13],c1[13]);
fa e15(a[14],b[14],c[14],s1[14],c1[14]);
fa e16(a[15],b[15],c[15],s1[15],c1[15]);

fa e17(a[16],b[16],c[16],s1[16],c1[16]);
fa e18(a[17],b[17],c[17],s1[17],c1[17]);
fa e19(a[18],b[18],c[18],s1[18],c1[18]);
fa e20(a[19],b[19],c[19],s1[19],c1[19]);
fa e21(a[20],b[20],c[20],s1[20],c1[20]);
fa e22(a[21],b[21],c[21],s1[21],c1[21]);
fa e23(a[22],b[22],c[22],s1[22],c1[22]);
fa e24(a[23],b[23],c[23],s1[23],c1[23]);

fa e25(a[24],b[24],c[24],s1[24],c1[24]);
fa e26(a[25],b[25],c[25],s1[25],c1[25]);
fa e27(a[26],b[26],c[26],s1[26],c1[26]);
fa e28(a[27],b[27],c[27],s1[27],c1[27]);
fa e29(a[28],b[28],c[28],s1[28],c1[28]);
fa e30(a[29],b[29],c[29],s1[29],c1[29]);
fa e31(a[30],b[30],c[30],s1[30],c1[30]);
fa e32(a[31],b[31],c[31],s1[31],c1[31]);

fa e33(a[32],b[32],c[32],s1[32],c1[32]);
fa e34(a[33],b[33],c[33],s1[33],c1[33]);
fa e35(a[34],b[34],c[34],s1[34],c1[34]);
fa e36(a[35],b[35],c[35],s1[35],c1[35]);
fa e37(a[36],b[36],c[36],s1[36],c1[36]);
fa e38(a[37],b[37],c[37],s1[37],c1[37]);
fa e39(a[38],b[38],c[38],s1[38],c1[38]);
fa e40(a[39],b[39],c[39],s1[39],c1[39]);

fa e41(a[40],b[40],c[40],s1[40],c1[40]); 
fa e42(a[41],b[41],c[41],s1[41],c1[41]);
fa e43(a[42],b[42],c[42],s1[42],c1[42]);
fa e44(a[43],b[43],c[43],s1[43],c1[43]);
fa e45(a[44],b[44],c[44],s1[44],c1[44]);
fa e46(a[45],b[45],c[45],s1[45],c1[45]);
fa e47(a[46],b[46],c[46],s1[46],c1[46]);
fa e48(a[47],b[47],c[47],s1[47],c1[47]);

fa e49(a[48],b[48],c[48],s1[48],c1[48]); 
fa e50(a[49],b[49],c[49],s1[49],c1[49]);
fa e51(a[50],b[50],c[50],s1[50],c1[50]);
fa e52(a[51],b[51],c[51],s1[51],c1[51]);
fa e53(a[52],b[52],c[52],s1[52],c1[52]);
fa e54(a[53],b[53],c[53],s1[53],c1[53]);
fa e55(a[54],b[54],c[54],s1[54],c1[54]);
fa e56(a[55],b[55],c[55],s1[55],c1[55]);

fa e57(a[56],b[56],c[56],s1[56],c1[56]); 
fa e58(a[57],b[57],c[57],s1[57],c1[57]);
fa e59(a[58],b[58],c[58],s1[58],c1[58]);
fa e60(a[59],b[59],c[59],s1[59],c1[59]);
fa e61(a[60],b[60],c[60],s1[60],c1[60]);
fa e62(a[61],b[61],c[61],s1[61],c1[61]);
fa e63(a[62],b[62],c[62],s1[62],c1[62]);
fa e64(a[63],b[63],c[63],s1[63],c1[63]);

assign s[0] =s1[0];

rca_64 r1({0,s1[63:1]},c1[63:0],s[64:1],0,cout);

endmodule
