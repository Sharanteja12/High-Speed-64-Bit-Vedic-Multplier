module csa_16 (a,b,c,s,cout);

input [15:0]a,b,c;
output [16:0] s;
output cout ;

wire [15:0] s1,c1;

fa e1(a[0],b[0],c[0],s1[0],c1[0]);
fa e2(a[1],b[1],c[1],s1[1],c1[1]);
fa e3(a[2],b[2],c[2],s1[2],c1[2]);
fa e4(a[3],b[3],c[3],s1[3],c1[3]);
fa e5(a[4],b[4],c[4],s1[4],c1[4]);
fa e6(a[5],b[5],c[5],s1[5],c1[5]);
fa e7(a[6],b[6],c[6],s1[6],c1[6]);
fa e8(a[7],b[7],c[7],s1[7],c1[7]);

fa e9(a[8],b[8],c[8],s1[8],c1[8]);
fa e10(a[9],b[9],c[9],s1[9],c1[9]);
fa e11(a[10],b[10],c[10],s1[10],c1[10]);
fa e12(a[11],b[11],c[11],s1[11],c1[11]);
fa e13(a[12],b[12],c[12],s1[12],c1[12]);
fa e14(a[13],b[13],c[13],s1[13],c1[13]);
fa e15(a[14],b[14],c[14],s1[14],c1[14]);
fa e16(a[15],b[15],c[15],s1[15],c1[15]);
assign s[0] =s1[0];

rca_16 r1({0,s1[15:1]},c1[15:0],s[16:1],0,cout);
endmodule
